`timescale 1ns/1ps
/*
    author : lbw
*/
module led_top(
    input   crtl,
    input   [31:0] num,
    output  LED0_CG,
    output  LED0_CF,
    output  LED0_CA,
    output  LED0_CB,
    output  LED0_CE,
    output  LED0_CD,
    output  LED0_CC,
    output  LED0_DP,
    output  DN0_K1,
    output  DN0_K2,
    output  DN0_K3,
    output  DN0_K4,
    output  LED1_CG,
    output  LED1_CF,
    output  LED1_CA,
    output  LED1_CB,
    output  LED1_CE,
    output  LED1_CD,
    output  LED1_CC,
    output  LED1_DP,
    output  DN1_K1,
    output  DN1_K2,
    output  DN1_K3,
    output  DN1_K4
);

    always @(*) begin
        
    end




endmodule