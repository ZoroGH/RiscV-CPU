`define I_BEQ  1
`define I_BNE  2
`define I_BLT  3
`define I_LW  4
`define I_SW  5
`define I_JAL  6
`define I_ADDI  7
`define I_ADD  8
`define I_SUB 9
`define I_MUL 10
`define I_MULH 11
`define I_BGE 12
`define I_XOR 13
`define I_AND 14
`define I_OR 15
`define I_LUI 16
`define I_AUIPC 17
`define I_ERR  5'd31
`define I_NULL 0