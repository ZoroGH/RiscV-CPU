`define I_BEQ  5'd1
`define I_BNE  5'd2
`define I_BLT  5'd3
`define I_LW  5'd4
`define I_SW  5'd5
`define I_JAL  5'd6
`define I_ADDI  5'd7
`define I_ADD  5'd8
`define I_SUB 5'd9
`define I_MUL 5'd10
`define I_MULH 5'd11
`define I_BGE 5'd12
`define I_XOR 5'd13
`define I_AND 5'd14
`define I_OR 5'd15
`define I_LUI 5'd16
`define I_AUIPC 5'd17
`define I_ERR  5'd31
`define I_NULL 5'd0
`define I_NOP 32'b00000000000000000000000000010011
`define I_ZEROS 32'd0
`define I_ONES 32'hFFFFFFFF