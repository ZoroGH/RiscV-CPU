module cpu_top(
    input clk
);

endmodule